entity vga_test is
end vga_test;

architecture vga_test of vga_test is
begin
end vga_test;
