entity vga is
end vga;

architecture vga of vga is
begin
end vga;
