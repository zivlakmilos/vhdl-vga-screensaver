entity main is
end main;

architecture main of main is
begin
end main;
